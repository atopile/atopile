* TPS54560 Peak Current-Mode Buck Converter Test
* 12V in, ~5V out, 5A load, 600kHz switching
* Uses the same TPS54560_TRANS model as the atopile design
*
.include models/TPS54560_TRANS.lib
*
* === Main circuit ===
V1 buck_vin 0 PULSE(0 12 0 10u 10u 10 10)
X1 boot comp buck_vin 0 sw rt buck_vin fb TPS54560_TRANS FS=600k
C_boot boot sw 100n
R_rt rt 0 162k
C_in buck_vin 0 30u
L1 sw power_out_hv 5.6u
C_out power_out_hv 0 88u
R_load power_out_hv 0 1
* Compensation network (TPS54560 reference design values)
R_comp comp comp_z 23.7k
C_comp1 comp_z 0 4.3n
C_comp2 comp 0 8.2p
* Feedback divider (Vout = 0.8 * (52.3k+10k)/10k = 4.984V)
R_top power_out_hv fb 52.3k
R_bottom fb 0 10k
*
.options reltol=0.003 abstol=1e-10 vntol=1e-5 gmin=1e-10 itl1=500 itl4=500 method=gear
.control
tran 200n 10m uic
wrdata /tmp/tps54560_test.txt v(power_out_hv) v(fb) i(L1) v(comp)
quit
.endc
.end
